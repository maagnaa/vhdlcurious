library IEEE;
use IEEE.std_logic_1164.all;

entity mux4_tb is
end entity mux4_tb;


architecture tb of mux4_tb is

 begin

end architecture tb;
