library IEEE;
use IEEE.std_logic_1164.all;

-- Why is the tb entity empty?!
entity mux2_tb is
end entity mux2_tb;


-- What are the steps we need to perform, which a testbench make?
-- 1. We need to instantiate a Device Under Test (DUT)...
-- 2. We need to apply some stimulus
-- 3. We need to confirm that the DUT behaves as we expect (aka. check the results)
-- (Hint! Look back at the testbench we used in smol_drill for ideas...)

architecture tb of mux2_tb is

 begin

end architecture tb;
