library IEEE; 
use IEEE.std_logic_1164.all;

entity mux4 is
  port(
    -- Oh dear... it sure is empty here.
  );
end;

architecture RTL of mux4 is

begin

end;
